module spi_clk_gen(  
    input wire clk,   
    input wire csn,    
    output reg sck       
);  
    // Frequency division coefficient parameter, SPI clock = clk / (2 * CLK_DIV)  
    parameter CLK_DIV = 4;  

    // Frequency counter that automatically switches the SCK level based on CLK_DIV  
    reg [15:0] clk_div_cnt = 16'd0;  

    always @(posedge clk or posedge csn) begin  
        if (csn) begin  
            clk_div_cnt <= 16'd0;  
            sck <= 1'b0;  
        end else begin  
            if (clk_div_cnt == (CLK_DIV - 1)) begin  
                clk_div_cnt <= 16'd0;  
                sck <= ~sck;  // Flip the clock  
            end else begin  
                clk_div_cnt <= clk_div_cnt + 16'd1;  
            end  
        end  
    end  
endmodule  

//https://www.chipverify.com/verilog/verilog-single-port-ram   
module single_port_sync_ram_master  
  # (parameter ADDR_WIDTH = 5,  
     parameter DATA_WIDTH = 24,  
     parameter DEPTH = 32  
    )  

  ( 	input 					clk,  
   		input [ADDR_WIDTH-1:0]	addr,  
   		inout [DATA_WIDTH-1:0]	data,  
   		input 					cs,  
   		input 					we,  
   		input 					oe  
  );  

  reg [DATA_WIDTH-1:0] 	tmp_data;  
  reg [DATA_WIDTH-1:0] 	mem [DEPTH];  

  always @ (posedge clk) begin  
    if (cs & we)  
      mem[addr] <= data;  
  end  

  always @ (posedge clk) begin  
    if (cs & !we)  
    	tmp_data <= mem[addr];  
  end  

  assign data = cs & oe & !we ? tmp_data : 'hz;   

  // Initialize RAM content  
  initial begin  
    // Initialize data at address 0.   
    mem[0] = 24'hABCDEF; // Example data  
    // Initialize other addresses to 0.  
    for (int i = 1; i < DEPTH; i = i + 1) begin  
      mem[i] = 24'h000000;  
    end  
  end  
  
endmodule  


module spi_master_top(  
    input wire clk,  
    input wire rstn,  
    output wire sck,     // Clock to slave  
    output reg csn,      // Chip select signal, active low  
    output reg mo,       // MOSI  
    input wire mi        // MISO  
);  

    // Parameter definition  
    parameter CLK_DIV = 4;  // SPI clock division ratio  

    // Internal registers  
    // reg [31:0] shift_reg;    
    reg [23:0] data_reg;    // 24-bit register to store data bits  
    reg [7:0] crc_reg;      // 8-bit register to store CRC checksum  
    reg [5:0] bit_cnt;      // Bit counter (0~31)  
    reg sck_en;             // SPI clock enable signal  
    reg time_cnt;           // Run count  

    // RAM control signals  
    reg [4:0] ram_addr;     
    reg ram_cs;              
    reg ram_we;              
    reg ram_oe;             
    wire [23:0] ram_data;    

    // State machine definition  
    typedef enum reg [2:0] {  
        IDLE,     // Idle state  
        WAIT,     // Waiting for RAM  
        WAIT2,  
        START,    // Start communication  
        TRANSFER  // Data transfer  
    } state_t;  
    state_t state;  

    // SPI clock signal connection  
    wire spi_sck;  
    
    // Instantiate the independent SPI clock generation module  
    spi_clk_gen #(  
        .CLK_DIV(CLK_DIV)  
    ) spi_clk_inst (  
        .clk(clk),  
        .csn(csn),  
        .sck(spi_sck)  
    );  
    
    // Connect the spi_sck signal generated by spi_clk_gen to the module's sck output  
    assign sck = spi_sck;   
    
    // CRC-8 SAE-J1850 polynomial  
    parameter CRC_POLY = 8'h1D;   

    // Instantiate RAM module  
    single_port_sync_ram_master #(  
        .ADDR_WIDTH(5),  
        .DATA_WIDTH(24),  
        .DEPTH(32)  
    ) ram_inst (  
        .clk(clk),  
        .addr(ram_addr),  
        .data(ram_data),  
        .cs(ram_cs),  
        .we(ram_we),  
        .oe(ram_oe)  
    );  

    // RAM Data Bus Driving Logic  
    assign ram_data = (ram_cs && ram_we) ? data_reg : 'hz;  
    
    reg [7:0] calculated_crc;  
    reg [23:0] temp_data;  
    integer i;   
    // Main logic for state machine  
    always @(posedge clk or negedge rstn) begin  
        if (!rstn) begin  
            csn <= 1'b1; // Chip select is disabled by default  
            data_reg <= 24'hA5A5A5; // Initialize data register   
            crc_reg <= 8'hFF;       // Initialize CRC register  
            bit_cnt <= 6'd0;  
            sck_en <= 1'b0;  
            state <= IDLE;  
            time_cnt <= 1'b1;  

        end else begin  
            case (state)  
                IDLE: begin  
                    csn <= 1'b1;    // Chip select inactive  
                    bit_cnt <= 6'd0;  
                    sck_en <= 1'b0;  
                    if (time_cnt > 1'b0) begin  
                        state <= WAIT;   

                    end else begin  
                        state <= IDLE;  
                    end  
                end  

                WAIT: begin  
                    // Read data from RAM into data_reg (upper half)  
                    ram_cs <= 1'b1;  
                    ram_we <= 1'b0;  
                    ram_oe <= 1'b1;  
                    ram_addr <= 5'd0;   

                    state <= WAIT2;  
                end  
                WAIT2: begin  
                    // Wait one clock cycle for ram_data to stabilize  
                    state <= START;  
                end   

                START: begin  
                    csn <= 1'b0;    // Pull chip select low to start communication  
                    sck_en <= 1'b1; // Enable SPI clock  
                    state <= TRANSFER;  
                    // Read data from RAM into data_reg (lower half)  
                    data_reg <= ram_data; // Load RAM data into data_reg  
                end  

                TRANSFER: begin  
                    if (bit_cnt == 6'd32) begin  // Transfer complete  
                        state <= IDLE;  
                        csn <= 1'b1;   // Disable chip select after transfer  
                        sck_en <= 1'b0;  // Disable SPI clock  
                        time_cnt <= time_cnt - 1'b1;  

                        /* Check CRC */  
                        // Recalculate CRC  
                        calculated_crc = 8'hFF;  // Initialize CRC  
                        temp_data = data_reg;    // Get current data  
                        for (i = 0; i < 24; i = i + 1) begin  
                            if (calculated_crc[7] ^ temp_data[23]) begin  
                                calculated_crc = (calculated_crc << 1) ^ CRC_POLY;  
                            end else begin  
                                calculated_crc = (calculated_crc << 1);  
                            end  
                            temp_data = temp_data << 1;  // Left shift data  
                        end  

                        // Compare recalculated CRC with received CRC  
                        if (calculated_crc != crc_reg) begin  
                            $display("CRC Error: Calculated CRC = %h, Received CRC = %h", calculated_crc, crc_reg);  
                        end else begin  
                            $display("CRC Check Passed");  
                        end  

                        // Write data_reg back to RAM  
                        // The assign statement already exists: ram_data = (ram_cs && ram_we) ? data_reg : 'hz; so only read/write permissions need to be changed  
                        ram_cs <= 1'b1;  
                        ram_we <= 1'b1;  
                        ram_oe <= 1'b0;  
                        ram_addr <= 5'd0; // Write address  
                    end  
                end  

                default: state <= IDLE;  
            endcase  
        end  
    end  

    // Handle data output on SCK rising edge  
    always @(posedge spi_sck or negedge rstn) begin  
        if (!rstn) begin  
            mo <= 1'b0;  
            crc_reg <= 8'hFF; // Initialize CRC register  
        end else if (!csn && sck_en) begin  
            if (bit_cnt < 24) begin  
                // Send data on SCK rising edge  
                mo <= data_reg[23];  
                // Dynamically update CRC register  
                if (crc_reg[7] ^ data_reg[23]) begin  // XOR operation  
                    crc_reg <= (crc_reg << 1) ^ CRC_POLY;  
                end else begin  
                    crc_reg <= (crc_reg << 1);  
                end  
            end else begin  
                // Send CRC checksum  
                mo <= crc_reg[7];  
            end  
        end  
    end  

    // Handle data reception on SCK falling edge  
    always @(negedge spi_sck or negedge rstn) begin  
        if (!rstn) begin  
            data_reg <= 24'hFFFFFF; // Initialize data register    
            bit_cnt <= 6'd0;  
        end else if (!csn && sck_en) begin  
            // Receive data on SCK falling edge  
            if (bit_cnt < 24) begin  
                data_reg  <= {data_reg [22:0], mi};  
            end else begin  
                // Receive CRC checksum  
                crc_reg <= {crc_reg[6:0], mi};  
            end   
            bit_cnt <= bit_cnt + 1'b1;  
        end  
    end  
endmodule